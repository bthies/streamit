//**********************************************************************
// Interface for input generator
//----------------------------------------------------------------------
//
//
//

package IInputGen;

import H264Types::*;
import GetPut::*;

interface IInputGen;

  // Interface for inter-module io
  interface Get#(InputGenOT) ioout;

endinterface

endpackage

